module buffer (B, A);
    input A;
    output B;

    assign B = A;


endmodule